.SUBCKT Transfer8_1 In_0 In_1 In_10 In_11 In_12 In_13 In_14 In_15 In_16 In_17 In_18 In_19 In_2 In_20 In_21 In_22 In_23 In_3 In_4 In_5 In_6 In_7 In_8 In_9 VDD VSS Y_0 Y_1 Y_10 Y_11 Y_12 Y_13 Y_14 Y_15 Y_2 Y_3 Y_4 Y_5 Y_6 Y_7 Y_8 Y_9
T1 T0_D In_2 VDD VSS nmos w=54.0n l=20n nfin=2 
T3 T2_D In_18 T0_D VSS nmos w=54.0n l=20n nfin=2 
T5 T4_D In_18 VDD VSS nmos w=54.0n l=20n nfin=2 
T7 T6_D In_20 T2_D VSS nmos w=54.0n l=20n nfin=2 
T9 T8_D In_20 T4_D VSS nmos w=54.0n l=20n nfin=2 
T11 T10_D In_20 VDD VSS nmos w=54.0n l=20n nfin=2 
T13 T12_D In_17 T6_D VSS nmos w=54.0n l=20n nfin=2 
T15 T14_D In_17 VDD VSS nmos w=54.0n l=20n nfin=2 
T17 T16_D In_17 T8_D VSS nmos w=54.0n l=20n nfin=2 
T19 T18_D In_17 T10_D VSS nmos w=54.0n l=20n nfin=2 
T21 T20_D In_16 T12_D VSS nmos w=54.0n l=20n nfin=2 
T23 T22_D In_16 VDD VSS nmos w=54.0n l=20n nfin=2 
T25 T24_D In_16 T14_D VSS nmos w=54.0n l=20n nfin=2 
T27 T26_D In_16 T16_D VSS nmos w=54.0n l=20n nfin=2 
T29 T28_D In_16 T18_D VSS nmos w=54.0n l=20n nfin=2 
T31 T30_D In_22 VDD VSS nmos w=54.0n l=20n nfin=2 
T33 T32_D In_22 T20_D VSS nmos w=54.0n l=20n nfin=2 
T35 T34_D In_22 T22_D VSS nmos w=54.0n l=20n nfin=2 
T37 T36_D In_22 T24_D VSS nmos w=54.0n l=20n nfin=2 
T39 T38_D In_22 T26_D VSS nmos w=54.0n l=20n nfin=2 
T41 T40_D In_22 T28_D VSS nmos w=54.0n l=20n nfin=2 
T43 T42_D In_23 T30_D VSS nmos w=54.0n l=20n nfin=2 
T45 T44_D In_23 VDD VSS nmos w=54.0n l=20n nfin=2 
T47 T46_D In_23 T32_D VSS nmos w=54.0n l=20n nfin=2 
T49 T48_D In_23 T34_D VSS nmos w=54.0n l=20n nfin=2 
T51 T50_D In_23 T36_D VSS nmos w=54.0n l=20n nfin=2 
T53 T52_D In_23 T38_D VSS nmos w=54.0n l=20n nfin=2 
T55 T54_D In_23 T40_D VSS nmos w=54.0n l=20n nfin=2 
T57 T56_D In_21 T42_D VSS nmos w=54.0n l=20n nfin=2 
T59 T58_D In_21 T44_D VSS nmos w=54.0n l=20n nfin=2 
T61 T60_D In_21 T46_D VSS nmos w=54.0n l=20n nfin=2 
T63 T62_D In_21 T48_D VSS nmos w=54.0n l=20n nfin=2 
T65 T64_D In_21 T50_D VSS nmos w=54.0n l=20n nfin=2 
T67 T66_D In_21 T52_D VSS nmos w=54.0n l=20n nfin=2 
T69 T68_D In_21 T54_D VSS nmos w=54.0n l=20n nfin=2 
T71 T70_D In_21 VDD VSS nmos w=54.0n l=20n nfin=2 
T73 T72_D In_15 T56_D VSS nmos w=54.0n l=20n nfin=2 
T75 T74_D In_15 T58_D VSS nmos w=54.0n l=20n nfin=2 
T77 T76_D In_15 VDD VSS nmos w=54.0n l=20n nfin=2 
T79 T78_D In_15 T60_D VSS nmos w=54.0n l=20n nfin=2 
T81 T80_D In_15 T62_D VSS nmos w=54.0n l=20n nfin=2 
T83 T82_D In_15 T64_D VSS nmos w=54.0n l=20n nfin=2 
T85 T84_D In_15 T66_D VSS nmos w=54.0n l=20n nfin=2 
T87 T86_D In_15 T68_D VSS nmos w=54.0n l=20n nfin=2 
T89 T88_D In_15 T70_D VSS nmos w=54.0n l=20n nfin=2 
T91 T90_D In_6 T72_D VSS nmos w=54.0n l=20n nfin=2 
T93 T92_D In_6 T74_D VSS nmos w=54.0n l=20n nfin=2 
T95 T94_D In_6 T76_D VSS nmos w=54.0n l=20n nfin=2 
T97 T96_D In_6 T78_D VSS nmos w=54.0n l=20n nfin=2 
T99 T98_D In_6 T80_D VSS nmos w=54.0n l=20n nfin=2 
T101 T100_D In_6 T82_D VSS nmos w=54.0n l=20n nfin=2 
T103 T102_D In_6 T84_D VSS nmos w=54.0n l=20n nfin=2 
T105 T104_D In_6 VDD VSS nmos w=54.0n l=20n nfin=2 
T107 T106_D In_6 T86_D VSS nmos w=54.0n l=20n nfin=2 
T109 T108_D In_6 T88_D VSS nmos w=54.0n l=20n nfin=2 
T111 T110_D In_19 T90_D VSS nmos w=54.0n l=20n nfin=2 
T113 T112_D In_19 T92_D VSS nmos w=54.0n l=20n nfin=2 
T115 T114_D In_19 T94_D VSS nmos w=54.0n l=20n nfin=2 
T117 T116_D In_19 T96_D VSS nmos w=54.0n l=20n nfin=2 
T119 T118_D In_19 T98_D VSS nmos w=54.0n l=20n nfin=2 
T121 T120_D In_19 T100_D VSS nmos w=54.0n l=20n nfin=2 
T123 T122_D In_19 T102_D VSS nmos w=54.0n l=20n nfin=2 
T125 T124_D In_19 VDD VSS nmos w=54.0n l=20n nfin=2 
T127 T126_D In_19 T104_D VSS nmos w=54.0n l=20n nfin=2 
T129 T128_D In_19 T106_D VSS nmos w=54.0n l=20n nfin=2 
T131 T130_D In_19 T108_D VSS nmos w=54.0n l=20n nfin=2 
T133 T132_D In_5 T110_D VSS nmos w=54.0n l=20n nfin=2 
T135 T134_D In_5 T112_D VSS nmos w=54.0n l=20n nfin=2 
T137 T136_D In_5 T114_D VSS nmos w=54.0n l=20n nfin=2 
T139 T138_D In_5 T116_D VSS nmos w=54.0n l=20n nfin=2 
T141 T140_D In_5 T118_D VSS nmos w=54.0n l=20n nfin=2 
T143 T142_D In_5 T120_D VSS nmos w=54.0n l=20n nfin=2 
T145 T144_D In_5 T122_D VSS nmos w=54.0n l=20n nfin=2 
T147 T146_D In_5 VDD VSS nmos w=54.0n l=20n nfin=2 
T149 T148_D In_5 T124_D VSS nmos w=54.0n l=20n nfin=2 
T151 T150_D In_5 T126_D VSS nmos w=54.0n l=20n nfin=2 
T153 T152_D In_5 T128_D VSS nmos w=54.0n l=20n nfin=2 
T155 T154_D In_5 T130_D VSS nmos w=54.0n l=20n nfin=2 
T157 T156_D In_4 T132_D VSS nmos w=54.0n l=20n nfin=2 
T159 T158_D In_4 T134_D VSS nmos w=54.0n l=20n nfin=2 
T161 T160_D In_4 T136_D VSS nmos w=54.0n l=20n nfin=2 
T163 T162_D In_4 T138_D VSS nmos w=54.0n l=20n nfin=2 
T165 T164_D In_4 T140_D VSS nmos w=54.0n l=20n nfin=2 
T167 T166_D In_4 T142_D VSS nmos w=54.0n l=20n nfin=2 
T169 T168_D In_4 VDD VSS nmos w=54.0n l=20n nfin=2 
T171 T170_D In_4 T144_D VSS nmos w=54.0n l=20n nfin=2 
T173 T172_D In_4 T146_D VSS nmos w=54.0n l=20n nfin=2 
T175 T174_D In_4 T148_D VSS nmos w=54.0n l=20n nfin=2 
T177 T176_D In_4 T150_D VSS nmos w=54.0n l=20n nfin=2 
T179 T178_D In_4 T152_D VSS nmos w=54.0n l=20n nfin=2 
T181 T180_D In_4 T154_D VSS nmos w=54.0n l=20n nfin=2 
T183 T182_D In_9 T156_D VSS nmos w=54.0n l=20n nfin=2 
T185 T184_D In_9 T158_D VSS nmos w=54.0n l=20n nfin=2 
T187 T186_D In_9 T160_D VSS nmos w=54.0n l=20n nfin=2 
T189 T188_D In_9 T162_D VSS nmos w=54.0n l=20n nfin=2 
T191 T190_D In_9 T164_D VSS nmos w=54.0n l=20n nfin=2 
T193 T192_D In_9 T166_D VSS nmos w=54.0n l=20n nfin=2 
T195 T194_D In_9 T168_D VSS nmos w=54.0n l=20n nfin=2 
T197 T196_D In_9 T170_D VSS nmos w=54.0n l=20n nfin=2 
T199 T198_D In_9 T172_D VSS nmos w=54.0n l=20n nfin=2 
T201 T200_D In_9 T174_D VSS nmos w=54.0n l=20n nfin=2 
T203 T202_D In_9 T176_D VSS nmos w=54.0n l=20n nfin=2 
T205 T204_D In_9 T178_D VSS nmos w=54.0n l=20n nfin=2 
T207 T206_D In_9 T180_D VSS nmos w=54.0n l=20n nfin=2 
T209 T208_D In_9 VDD VSS nmos w=54.0n l=20n nfin=2 
T211 T210_D In_8 T182_D VSS nmos w=54.0n l=20n nfin=2 
T213 T212_D In_8 T184_D VSS nmos w=54.0n l=20n nfin=2 
T215 T214_D In_8 T186_D VSS nmos w=54.0n l=20n nfin=2 
T217 T216_D In_8 T188_D VSS nmos w=54.0n l=20n nfin=2 
T219 T218_D In_8 T190_D VSS nmos w=54.0n l=20n nfin=2 
T221 T220_D In_8 T192_D VSS nmos w=54.0n l=20n nfin=2 
T223 T222_D In_8 T194_D VSS nmos w=54.0n l=20n nfin=2 
T225 T224_D In_8 T196_D VSS nmos w=54.0n l=20n nfin=2 
T227 T226_D In_8 T198_D VSS nmos w=54.0n l=20n nfin=2 
T229 T228_D In_8 T200_D VSS nmos w=54.0n l=20n nfin=2 
T231 T230_D In_8 T202_D VSS nmos w=54.0n l=20n nfin=2 
T233 T232_D In_8 T204_D VSS nmos w=54.0n l=20n nfin=2 
T235 T234_D In_8 T206_D VSS nmos w=54.0n l=20n nfin=2 
T237 T236_D In_8 VDD VSS nmos w=54.0n l=20n nfin=2 
T239 T238_D In_8 T208_D VSS nmos w=54.0n l=20n nfin=2 
T241 T240_D In_7 T210_D VSS nmos w=54.0n l=20n nfin=2 
T243 T242_D In_7 T212_D VSS nmos w=54.0n l=20n nfin=2 
T245 T244_D In_7 T214_D VSS nmos w=54.0n l=20n nfin=2 
T247 T246_D In_7 T216_D VSS nmos w=54.0n l=20n nfin=2 
T249 T248_D In_7 T218_D VSS nmos w=54.0n l=20n nfin=2 
T251 T250_D In_7 T220_D VSS nmos w=54.0n l=20n nfin=2 
T253 T252_D In_7 T222_D VSS nmos w=54.0n l=20n nfin=2 
T255 T254_D In_7 T224_D VSS nmos w=54.0n l=20n nfin=2 
T257 T256_D In_7 T226_D VSS nmos w=54.0n l=20n nfin=2 
T259 T258_D In_7 T228_D VSS nmos w=54.0n l=20n nfin=2 
T261 T260_D In_7 T230_D VSS nmos w=54.0n l=20n nfin=2 
T263 T262_D In_7 T232_D VSS nmos w=54.0n l=20n nfin=2 
T265 T264_D In_7 VDD VSS nmos w=54.0n l=20n nfin=2 
T267 T266_D In_7 T234_D VSS nmos w=54.0n l=20n nfin=2 
T269 T268_D In_7 T236_D VSS nmos w=54.0n l=20n nfin=2 
T271 T270_D In_7 T238_D VSS nmos w=54.0n l=20n nfin=2 
T273 T272_D In_3 T240_D VSS nmos w=54.0n l=20n nfin=2 
T275 T274_D In_3 T242_D VSS nmos w=54.0n l=20n nfin=2 
T277 T276_D In_3 T244_D VSS nmos w=54.0n l=20n nfin=2 
T279 T278_D In_3 T246_D VSS nmos w=54.0n l=20n nfin=2 
T281 T280_D In_3 T248_D VSS nmos w=54.0n l=20n nfin=2 
T283 T282_D In_3 VDD VSS nmos w=54.0n l=20n nfin=2 
T285 T284_D In_3 T250_D VSS nmos w=54.0n l=20n nfin=2 
T287 T286_D In_3 T252_D VSS nmos w=54.0n l=20n nfin=2 
T289 T288_D In_3 T254_D VSS nmos w=54.0n l=20n nfin=2 
T291 T290_D In_3 T256_D VSS nmos w=54.0n l=20n nfin=2 
T293 T292_D In_3 T258_D VSS nmos w=54.0n l=20n nfin=2 
T295 T294_D In_3 T260_D VSS nmos w=54.0n l=20n nfin=2 
T297 T296_D In_3 T262_D VSS nmos w=54.0n l=20n nfin=2 
T299 T298_D In_3 T264_D VSS nmos w=54.0n l=20n nfin=2 
T301 T300_D In_3 T266_D VSS nmos w=54.0n l=20n nfin=2 
T303 T302_D In_3 T268_D VSS nmos w=54.0n l=20n nfin=2 
T305 T304_D In_3 T270_D VSS nmos w=54.0n l=20n nfin=2 
T307 T306_D In_13 T272_D VSS nmos w=54.0n l=20n nfin=2 
T309 T308_D In_13 T274_D VSS nmos w=54.0n l=20n nfin=2 
T311 T310_D In_13 VDD VSS nmos w=54.0n l=20n nfin=2 
T313 T312_D In_13 T276_D VSS nmos w=54.0n l=20n nfin=2 
T315 T314_D In_13 VSS VSS nmos w=54.0n l=20n nfin=2 
T317 T316_D In_13 T280_D VSS nmos w=54.0n l=20n nfin=2 
T319 T318_D In_13 T276_D VSS nmos w=54.0n l=20n nfin=2 
T321 T320_D In_13 T284_D VSS nmos w=54.0n l=20n nfin=2 
T323 T322_D In_13 T280_D VSS nmos w=54.0n l=20n nfin=2 
T325 T324_D In_13 T288_D VSS nmos w=54.0n l=20n nfin=2 
T327 T326_D In_13 T284_D VSS nmos w=54.0n l=20n nfin=2 
T329 T328_D In_13 T292_D VSS nmos w=54.0n l=20n nfin=2 
T331 T330_D In_13 T288_D VSS nmos w=54.0n l=20n nfin=2 
T333 T332_D In_13 T296_D VSS nmos w=54.0n l=20n nfin=2 
T335 T334_D In_13 T292_D VSS nmos w=54.0n l=20n nfin=2 
T337 T336_D In_13 T300_D VSS nmos w=54.0n l=20n nfin=2 
T339 T338_D In_13 T296_D VSS nmos w=54.0n l=20n nfin=2 
T341 T340_D In_13 T300_D VSS nmos w=54.0n l=20n nfin=2 
T343 T342_D In_14 T306_D VSS nmos w=54.0n l=20n nfin=2 
T345 T344_D In_14 T308_D VSS nmos w=54.0n l=20n nfin=2 
T347 T346_D In_14 T310_D VSS nmos w=54.0n l=20n nfin=2 
T349 T348_D In_14 VDD VSS nmos w=54.0n l=20n nfin=2 
T351 T350_D In_14 T310_D VSS nmos w=54.0n l=20n nfin=2 
T353 T352_D In_14 T312_D VSS nmos w=54.0n l=20n nfin=2 
T355 T354_D In_14 VSS VSS nmos w=54.0n l=20n nfin=2 
T357 T356_D In_14 T316_D VSS nmos w=54.0n l=20n nfin=2 
T359 T358_D In_14 T312_D VSS nmos w=54.0n l=20n nfin=2 
T361 T360_D In_14 T320_D VSS nmos w=54.0n l=20n nfin=2 
T363 T362_D In_14 T316_D VSS nmos w=54.0n l=20n nfin=2 
T365 T364_D In_14 T324_D VSS nmos w=54.0n l=20n nfin=2 
T367 T366_D In_14 T320_D VSS nmos w=54.0n l=20n nfin=2 
T369 T368_D In_14 T328_D VSS nmos w=54.0n l=20n nfin=2 
T371 T370_D In_14 T324_D VSS nmos w=54.0n l=20n nfin=2 
T373 T372_D In_14 T332_D VSS nmos w=54.0n l=20n nfin=2 
T375 T374_D In_14 T328_D VSS nmos w=54.0n l=20n nfin=2 
T377 T376_D In_14 T336_D VSS nmos w=54.0n l=20n nfin=2 
T379 T378_D In_14 T332_D VSS nmos w=54.0n l=20n nfin=2 
T381 T380_D In_14 T336_D VSS nmos w=54.0n l=20n nfin=2 
T383 T382_D In_14 VSS VSS nmos w=54.0n l=20n nfin=2 
T385 T384_D In_12 T342_D VSS nmos w=54.0n l=20n nfin=2 
T387 T386_D In_12 T344_D VSS nmos w=54.0n l=20n nfin=2 
T389 T388_D In_12 VSS VSS nmos w=54.0n l=20n nfin=2 
T391 T390_D In_12 T346_D VSS nmos w=54.0n l=20n nfin=2 
T393 T392_D In_12 T350_D VSS nmos w=54.0n l=20n nfin=2 
T395 T394_D In_12 T352_D VSS nmos w=54.0n l=20n nfin=2 
T397 T396_D In_12 VSS VSS nmos w=54.0n l=20n nfin=2 
T399 T398_D In_12 T356_D VSS nmos w=54.0n l=20n nfin=2 
T401 T400_D In_12 T352_D VSS nmos w=54.0n l=20n nfin=2 
T403 T402_D In_12 T360_D VSS nmos w=54.0n l=20n nfin=2 
T405 T404_D In_12 T356_D VSS nmos w=54.0n l=20n nfin=2 
T407 T406_D In_12 T364_D VSS nmos w=54.0n l=20n nfin=2 
T409 T408_D In_12 T360_D VSS nmos w=54.0n l=20n nfin=2 
T411 T410_D In_12 T368_D VSS nmos w=54.0n l=20n nfin=2 
T413 T412_D In_12 T364_D VSS nmos w=54.0n l=20n nfin=2 
T415 T414_D In_12 T372_D VSS nmos w=54.0n l=20n nfin=2 
T417 T416_D In_12 T368_D VSS nmos w=54.0n l=20n nfin=2 
T419 T418_D In_12 T376_D VSS nmos w=54.0n l=20n nfin=2 
T421 T420_D In_12 T372_D VSS nmos w=54.0n l=20n nfin=2 
T423 T422_D In_12 T376_D VSS nmos w=54.0n l=20n nfin=2 
T425 T424_D In_12 VSS VSS nmos w=54.0n l=20n nfin=2 
T427 T426_D In_10 T384_D VSS nmos w=54.0n l=20n nfin=2 
T429 T428_D In_10 T386_D VSS nmos w=54.0n l=20n nfin=2 
T431 T430_D In_10 T388_D VSS nmos w=54.0n l=20n nfin=2 
T433 T432_D In_10 T390_D VSS nmos w=54.0n l=20n nfin=2 
T435 T434_D In_10 T392_D VSS nmos w=54.0n l=20n nfin=2 
T437 T436_D In_10 T396_D VSS nmos w=54.0n l=20n nfin=2 
T439 T438_D In_10 T400_D VSS nmos w=54.0n l=20n nfin=2 
T441 T440_D In_10 T404_D VSS nmos w=54.0n l=20n nfin=2 
T443 T442_D In_10 T408_D VSS nmos w=54.0n l=20n nfin=2 
T445 T444_D In_10 T412_D VSS nmos w=54.0n l=20n nfin=2 
T447 T446_D In_10 T416_D VSS nmos w=54.0n l=20n nfin=2 
T449 T448_D In_10 T420_D VSS nmos w=54.0n l=20n nfin=2 
T451 T450_D In_10 T422_D VSS nmos w=54.0n l=20n nfin=2 
T453 T452_D In_10 T424_D VSS nmos w=54.0n l=20n nfin=2 
T455 T454_D In_11 T426_D VSS nmos w=54.0n l=20n nfin=2 
T457 T456_D In_11 T428_D VSS nmos w=54.0n l=20n nfin=2 
T459 T458_D In_11 VDD VSS nmos w=54.0n l=20n nfin=2 
T461 T460_D In_11 T430_D VSS nmos w=54.0n l=20n nfin=2 
T463 T462_D In_11 T432_D VSS nmos w=54.0n l=20n nfin=2 
T465 T464_D In_11 T434_D VSS nmos w=54.0n l=20n nfin=2 
T467 T466_D In_11 T436_D VSS nmos w=54.0n l=20n nfin=2 
T469 T468_D In_11 T438_D VSS nmos w=54.0n l=20n nfin=2 
T471 T470_D In_11 T440_D VSS nmos w=54.0n l=20n nfin=2 
T473 T472_D In_11 T442_D VSS nmos w=54.0n l=20n nfin=2 
T475 T474_D In_11 T444_D VSS nmos w=54.0n l=20n nfin=2 
T477 T476_D In_11 T446_D VSS nmos w=54.0n l=20n nfin=2 
T479 T478_D In_11 T448_D VSS nmos w=54.0n l=20n nfin=2 
T481 T480_D In_11 T450_D VSS nmos w=54.0n l=20n nfin=2 
T483 T482_D In_11 T452_D VSS nmos w=54.0n l=20n nfin=2 
T485 Y_0 In_1 T454_D VSS nmos w=54.0n l=20n nfin=2 
T487 Y_1 In_1 T456_D VSS nmos w=54.0n l=20n nfin=2 
T489 Y_2 In_1 T458_D VSS nmos w=54.0n l=20n nfin=2 
T491 Y_3 In_1 VDD VSS nmos w=54.0n l=20n nfin=2 
T493 Y_4 In_1 T460_D VSS nmos w=54.0n l=20n nfin=2 
T495 Y_5 In_1 T462_D VSS nmos w=54.0n l=20n nfin=2 
T497 Y_6 In_1 T464_D VSS nmos w=54.0n l=20n nfin=2 
T499 Y_7 In_1 T466_D VSS nmos w=54.0n l=20n nfin=2 
T501 Y_8 In_1 T468_D VSS nmos w=54.0n l=20n nfin=2 
T503 Y_9 In_1 T470_D VSS nmos w=54.0n l=20n nfin=2 
T505 Y_10 In_1 T472_D VSS nmos w=54.0n l=20n nfin=2 
T507 Y_11 In_1 T474_D VSS nmos w=54.0n l=20n nfin=2 
T509 Y_12 In_1 T476_D VSS nmos w=54.0n l=20n nfin=2 
T511 Y_13 In_1 T478_D VSS nmos w=54.0n l=20n nfin=2 
T513 Y_14 In_1 T480_D VSS nmos w=54.0n l=20n nfin=2 
T515 Y_15 In_1 T482_D VSS nmos w=54.0n l=20n nfin=2 
T0 T0_D In_2 VSS VDD pmos w=54.0n l=20n nfin=2 
T2 T2_D In_18 T0_D VDD pmos w=54.0n l=20n nfin=2 
T4 T4_D In_18 VSS VDD pmos w=54.0n l=20n nfin=2 
T6 T6_D In_20 T2_D VDD pmos w=54.0n l=20n nfin=2 
T8 T8_D In_20 T4_D VDD pmos w=54.0n l=20n nfin=2 
T10 T10_D In_20 VSS VDD pmos w=54.0n l=20n nfin=2 
T12 T12_D In_17 T6_D VDD pmos w=54.0n l=20n nfin=2 
T14 T14_D In_17 VSS VDD pmos w=54.0n l=20n nfin=2 
T16 T16_D In_17 T8_D VDD pmos w=54.0n l=20n nfin=2 
T18 T18_D In_17 T10_D VDD pmos w=54.0n l=20n nfin=2 
T20 T20_D In_16 T12_D VDD pmos w=54.0n l=20n nfin=2 
T22 T22_D In_16 VSS VDD pmos w=54.0n l=20n nfin=2 
T24 T24_D In_16 T14_D VDD pmos w=54.0n l=20n nfin=2 
T26 T26_D In_16 T16_D VDD pmos w=54.0n l=20n nfin=2 
T28 T28_D In_16 T18_D VDD pmos w=54.0n l=20n nfin=2 
T30 T30_D In_22 VSS VDD pmos w=54.0n l=20n nfin=2 
T32 T32_D In_22 T20_D VDD pmos w=54.0n l=20n nfin=2 
T34 T34_D In_22 T22_D VDD pmos w=54.0n l=20n nfin=2 
T36 T36_D In_22 T24_D VDD pmos w=54.0n l=20n nfin=2 
T38 T38_D In_22 T26_D VDD pmos w=54.0n l=20n nfin=2 
T40 T40_D In_22 T28_D VDD pmos w=54.0n l=20n nfin=2 
T42 T42_D In_23 T30_D VDD pmos w=54.0n l=20n nfin=2 
T44 T44_D In_23 VSS VDD pmos w=54.0n l=20n nfin=2 
T46 T46_D In_23 T32_D VDD pmos w=54.0n l=20n nfin=2 
T48 T48_D In_23 T34_D VDD pmos w=54.0n l=20n nfin=2 
T50 T50_D In_23 T36_D VDD pmos w=54.0n l=20n nfin=2 
T52 T52_D In_23 T38_D VDD pmos w=54.0n l=20n nfin=2 
T54 T54_D In_23 T40_D VDD pmos w=54.0n l=20n nfin=2 
T56 T56_D In_21 T42_D VDD pmos w=54.0n l=20n nfin=2 
T58 T58_D In_21 T44_D VDD pmos w=54.0n l=20n nfin=2 
T60 T60_D In_21 T46_D VDD pmos w=54.0n l=20n nfin=2 
T62 T62_D In_21 T48_D VDD pmos w=54.0n l=20n nfin=2 
T64 T64_D In_21 T50_D VDD pmos w=54.0n l=20n nfin=2 
T66 T66_D In_21 T52_D VDD pmos w=54.0n l=20n nfin=2 
T68 T68_D In_21 T54_D VDD pmos w=54.0n l=20n nfin=2 
T70 T70_D In_21 VSS VDD pmos w=54.0n l=20n nfin=2 
T72 T72_D In_15 T56_D VDD pmos w=54.0n l=20n nfin=2 
T74 T74_D In_15 T58_D VDD pmos w=54.0n l=20n nfin=2 
T76 T76_D In_15 VSS VDD pmos w=54.0n l=20n nfin=2 
T78 T78_D In_15 T60_D VDD pmos w=54.0n l=20n nfin=2 
T80 T80_D In_15 T62_D VDD pmos w=54.0n l=20n nfin=2 
T82 T82_D In_15 T64_D VDD pmos w=54.0n l=20n nfin=2 
T84 T84_D In_15 T66_D VDD pmos w=54.0n l=20n nfin=2 
T86 T86_D In_15 T68_D VDD pmos w=54.0n l=20n nfin=2 
T88 T88_D In_15 T70_D VDD pmos w=54.0n l=20n nfin=2 
T90 T90_D In_6 T72_D VDD pmos w=54.0n l=20n nfin=2 
T92 T92_D In_6 T74_D VDD pmos w=54.0n l=20n nfin=2 
T94 T94_D In_6 T76_D VDD pmos w=54.0n l=20n nfin=2 
T96 T96_D In_6 T78_D VDD pmos w=54.0n l=20n nfin=2 
T98 T98_D In_6 T80_D VDD pmos w=54.0n l=20n nfin=2 
T100 T100_D In_6 T82_D VDD pmos w=54.0n l=20n nfin=2 
T102 T102_D In_6 T84_D VDD pmos w=54.0n l=20n nfin=2 
T104 T104_D In_6 VSS VDD pmos w=54.0n l=20n nfin=2 
T106 T106_D In_6 T86_D VDD pmos w=54.0n l=20n nfin=2 
T108 T108_D In_6 T88_D VDD pmos w=54.0n l=20n nfin=2 
T110 T110_D In_19 T90_D VDD pmos w=54.0n l=20n nfin=2 
T112 T112_D In_19 T92_D VDD pmos w=54.0n l=20n nfin=2 
T114 T114_D In_19 T94_D VDD pmos w=54.0n l=20n nfin=2 
T116 T116_D In_19 T96_D VDD pmos w=54.0n l=20n nfin=2 
T118 T118_D In_19 T98_D VDD pmos w=54.0n l=20n nfin=2 
T120 T120_D In_19 T100_D VDD pmos w=54.0n l=20n nfin=2 
T122 T122_D In_19 T102_D VDD pmos w=54.0n l=20n nfin=2 
T124 T124_D In_19 VSS VDD pmos w=54.0n l=20n nfin=2 
T126 T126_D In_19 T104_D VDD pmos w=54.0n l=20n nfin=2 
T128 T128_D In_19 T106_D VDD pmos w=54.0n l=20n nfin=2 
T130 T130_D In_19 T108_D VDD pmos w=54.0n l=20n nfin=2 
T132 T132_D In_5 T110_D VDD pmos w=54.0n l=20n nfin=2 
T134 T134_D In_5 T112_D VDD pmos w=54.0n l=20n nfin=2 
T136 T136_D In_5 T114_D VDD pmos w=54.0n l=20n nfin=2 
T138 T138_D In_5 T116_D VDD pmos w=54.0n l=20n nfin=2 
T140 T140_D In_5 T118_D VDD pmos w=54.0n l=20n nfin=2 
T142 T142_D In_5 T120_D VDD pmos w=54.0n l=20n nfin=2 
T144 T144_D In_5 T122_D VDD pmos w=54.0n l=20n nfin=2 
T146 T146_D In_5 VSS VDD pmos w=54.0n l=20n nfin=2 
T148 T148_D In_5 T124_D VDD pmos w=54.0n l=20n nfin=2 
T150 T150_D In_5 T126_D VDD pmos w=54.0n l=20n nfin=2 
T152 T152_D In_5 T128_D VDD pmos w=54.0n l=20n nfin=2 
T154 T154_D In_5 T130_D VDD pmos w=54.0n l=20n nfin=2 
T156 T156_D In_4 T132_D VDD pmos w=54.0n l=20n nfin=2 
T158 T158_D In_4 T134_D VDD pmos w=54.0n l=20n nfin=2 
T160 T160_D In_4 T136_D VDD pmos w=54.0n l=20n nfin=2 
T162 T162_D In_4 T138_D VDD pmos w=54.0n l=20n nfin=2 
T164 T164_D In_4 T140_D VDD pmos w=54.0n l=20n nfin=2 
T166 T166_D In_4 T142_D VDD pmos w=54.0n l=20n nfin=2 
T168 T168_D In_4 VSS VDD pmos w=54.0n l=20n nfin=2 
T170 T170_D In_4 T144_D VDD pmos w=54.0n l=20n nfin=2 
T172 T172_D In_4 T146_D VDD pmos w=54.0n l=20n nfin=2 
T174 T174_D In_4 T148_D VDD pmos w=54.0n l=20n nfin=2 
T176 T176_D In_4 T150_D VDD pmos w=54.0n l=20n nfin=2 
T178 T178_D In_4 T152_D VDD pmos w=54.0n l=20n nfin=2 
T180 T180_D In_4 T154_D VDD pmos w=54.0n l=20n nfin=2 
T182 T182_D In_9 T156_D VDD pmos w=54.0n l=20n nfin=2 
T184 T184_D In_9 T158_D VDD pmos w=54.0n l=20n nfin=2 
T186 T186_D In_9 T160_D VDD pmos w=54.0n l=20n nfin=2 
T188 T188_D In_9 T162_D VDD pmos w=54.0n l=20n nfin=2 
T190 T190_D In_9 T164_D VDD pmos w=54.0n l=20n nfin=2 
T192 T192_D In_9 T166_D VDD pmos w=54.0n l=20n nfin=2 
T194 T194_D In_9 T168_D VDD pmos w=54.0n l=20n nfin=2 
T196 T196_D In_9 T170_D VDD pmos w=54.0n l=20n nfin=2 
T198 T198_D In_9 T172_D VDD pmos w=54.0n l=20n nfin=2 
T200 T200_D In_9 T174_D VDD pmos w=54.0n l=20n nfin=2 
T202 T202_D In_9 T176_D VDD pmos w=54.0n l=20n nfin=2 
T204 T204_D In_9 T178_D VDD pmos w=54.0n l=20n nfin=2 
T206 T206_D In_9 T180_D VDD pmos w=54.0n l=20n nfin=2 
T208 T208_D In_9 VSS VDD pmos w=54.0n l=20n nfin=2 
T210 T210_D In_8 T182_D VDD pmos w=54.0n l=20n nfin=2 
T212 T212_D In_8 T184_D VDD pmos w=54.0n l=20n nfin=2 
T214 T214_D In_8 T186_D VDD pmos w=54.0n l=20n nfin=2 
T216 T216_D In_8 T188_D VDD pmos w=54.0n l=20n nfin=2 
T218 T218_D In_8 T190_D VDD pmos w=54.0n l=20n nfin=2 
T220 T220_D In_8 T192_D VDD pmos w=54.0n l=20n nfin=2 
T222 T222_D In_8 T194_D VDD pmos w=54.0n l=20n nfin=2 
T224 T224_D In_8 T196_D VDD pmos w=54.0n l=20n nfin=2 
T226 T226_D In_8 T198_D VDD pmos w=54.0n l=20n nfin=2 
T228 T228_D In_8 T200_D VDD pmos w=54.0n l=20n nfin=2 
T230 T230_D In_8 T202_D VDD pmos w=54.0n l=20n nfin=2 
T232 T232_D In_8 T204_D VDD pmos w=54.0n l=20n nfin=2 
T234 T234_D In_8 T206_D VDD pmos w=54.0n l=20n nfin=2 
T236 T236_D In_8 VSS VDD pmos w=54.0n l=20n nfin=2 
T238 T238_D In_8 T208_D VDD pmos w=54.0n l=20n nfin=2 
T240 T240_D In_7 T210_D VDD pmos w=54.0n l=20n nfin=2 
T242 T242_D In_7 T212_D VDD pmos w=54.0n l=20n nfin=2 
T244 T244_D In_7 T214_D VDD pmos w=54.0n l=20n nfin=2 
T246 T246_D In_7 T216_D VDD pmos w=54.0n l=20n nfin=2 
T248 T248_D In_7 T218_D VDD pmos w=54.0n l=20n nfin=2 
T250 T250_D In_7 T220_D VDD pmos w=54.0n l=20n nfin=2 
T252 T252_D In_7 T222_D VDD pmos w=54.0n l=20n nfin=2 
T254 T254_D In_7 T224_D VDD pmos w=54.0n l=20n nfin=2 
T256 T256_D In_7 T226_D VDD pmos w=54.0n l=20n nfin=2 
T258 T258_D In_7 T228_D VDD pmos w=54.0n l=20n nfin=2 
T260 T260_D In_7 T230_D VDD pmos w=54.0n l=20n nfin=2 
T262 T262_D In_7 T232_D VDD pmos w=54.0n l=20n nfin=2 
T264 T264_D In_7 VSS VDD pmos w=54.0n l=20n nfin=2 
T266 T266_D In_7 T234_D VDD pmos w=54.0n l=20n nfin=2 
T268 T268_D In_7 T236_D VDD pmos w=54.0n l=20n nfin=2 
T270 T270_D In_7 T238_D VDD pmos w=54.0n l=20n nfin=2 
T272 T272_D In_3 T240_D VDD pmos w=54.0n l=20n nfin=2 
T274 T274_D In_3 T242_D VDD pmos w=54.0n l=20n nfin=2 
T276 T276_D In_3 T244_D VDD pmos w=54.0n l=20n nfin=2 
T278 T278_D In_3 T246_D VDD pmos w=54.0n l=20n nfin=2 
T280 T280_D In_3 T248_D VDD pmos w=54.0n l=20n nfin=2 
T282 T282_D In_3 VSS VDD pmos w=54.0n l=20n nfin=2 
T284 T284_D In_3 T250_D VDD pmos w=54.0n l=20n nfin=2 
T286 T286_D In_3 T252_D VDD pmos w=54.0n l=20n nfin=2 
T288 T288_D In_3 T254_D VDD pmos w=54.0n l=20n nfin=2 
T290 T290_D In_3 T256_D VDD pmos w=54.0n l=20n nfin=2 
T292 T292_D In_3 T258_D VDD pmos w=54.0n l=20n nfin=2 
T294 T294_D In_3 T260_D VDD pmos w=54.0n l=20n nfin=2 
T296 T296_D In_3 T262_D VDD pmos w=54.0n l=20n nfin=2 
T298 T298_D In_3 T264_D VDD pmos w=54.0n l=20n nfin=2 
T300 T300_D In_3 T266_D VDD pmos w=54.0n l=20n nfin=2 
T302 T302_D In_3 T268_D VDD pmos w=54.0n l=20n nfin=2 
T304 T304_D In_3 T270_D VDD pmos w=54.0n l=20n nfin=2 
T306 T306_D In_13 T272_D VDD pmos w=54.0n l=20n nfin=2 
T308 T308_D In_13 T274_D VDD pmos w=54.0n l=20n nfin=2 
T310 T310_D In_13 VSS VDD pmos w=54.0n l=20n nfin=2 
T312 T312_D In_13 T276_D VDD pmos w=54.0n l=20n nfin=2 
T314 T314_D In_13 T278_D VDD pmos w=54.0n l=20n nfin=2 
T316 T316_D In_13 T280_D VDD pmos w=54.0n l=20n nfin=2 
T318 T318_D In_13 T282_D VDD pmos w=54.0n l=20n nfin=2 
T320 T320_D In_13 T284_D VDD pmos w=54.0n l=20n nfin=2 
T322 T322_D In_13 T286_D VDD pmos w=54.0n l=20n nfin=2 
T324 T324_D In_13 T288_D VDD pmos w=54.0n l=20n nfin=2 
T326 T326_D In_13 T290_D VDD pmos w=54.0n l=20n nfin=2 
T328 T328_D In_13 T292_D VDD pmos w=54.0n l=20n nfin=2 
T330 T330_D In_13 T294_D VDD pmos w=54.0n l=20n nfin=2 
T332 T332_D In_13 T296_D VDD pmos w=54.0n l=20n nfin=2 
T334 T334_D In_13 T298_D VDD pmos w=54.0n l=20n nfin=2 
T336 T336_D In_13 T300_D VDD pmos w=54.0n l=20n nfin=2 
T338 T338_D In_13 T302_D VDD pmos w=54.0n l=20n nfin=2 
T340 T340_D In_13 T304_D VDD pmos w=54.0n l=20n nfin=2 
T342 T342_D In_14 T306_D VDD pmos w=54.0n l=20n nfin=2 
T344 T344_D In_14 T308_D VDD pmos w=54.0n l=20n nfin=2 
T346 T346_D In_14 T310_D VDD pmos w=54.0n l=20n nfin=2 
T348 T348_D In_14 VSS VDD pmos w=54.0n l=20n nfin=2 
T350 T350_D In_14 T310_D VDD pmos w=54.0n l=20n nfin=2 
T352 T352_D In_14 T312_D VDD pmos w=54.0n l=20n nfin=2 
T354 T354_D In_14 T314_D VDD pmos w=54.0n l=20n nfin=2 
T356 T356_D In_14 T316_D VDD pmos w=54.0n l=20n nfin=2 
T358 T358_D In_14 T318_D VDD pmos w=54.0n l=20n nfin=2 
T360 T360_D In_14 T320_D VDD pmos w=54.0n l=20n nfin=2 
T362 T362_D In_14 T322_D VDD pmos w=54.0n l=20n nfin=2 
T364 T364_D In_14 T324_D VDD pmos w=54.0n l=20n nfin=2 
T366 T366_D In_14 T326_D VDD pmos w=54.0n l=20n nfin=2 
T368 T368_D In_14 T328_D VDD pmos w=54.0n l=20n nfin=2 
T370 T370_D In_14 T330_D VDD pmos w=54.0n l=20n nfin=2 
T372 T372_D In_14 T332_D VDD pmos w=54.0n l=20n nfin=2 
T374 T374_D In_14 T334_D VDD pmos w=54.0n l=20n nfin=2 
T376 T376_D In_14 T336_D VDD pmos w=54.0n l=20n nfin=2 
T378 T378_D In_14 T338_D VDD pmos w=54.0n l=20n nfin=2 
T380 T380_D In_14 T340_D VDD pmos w=54.0n l=20n nfin=2 
T382 T382_D In_14 T310_D VDD pmos w=54.0n l=20n nfin=2 
T384 T384_D In_12 T342_D VDD pmos w=54.0n l=20n nfin=2 
T386 T386_D In_12 T344_D VDD pmos w=54.0n l=20n nfin=2 
T388 T388_D In_12 VDD VDD pmos w=54.0n l=20n nfin=2 
T390 T390_D In_12 T346_D VDD pmos w=54.0n l=20n nfin=2 
T392 T392_D In_12 T348_D VDD pmos w=54.0n l=20n nfin=2 
T394 T394_D In_12 T352_D VDD pmos w=54.0n l=20n nfin=2 
T396 T396_D In_12 T354_D VDD pmos w=54.0n l=20n nfin=2 
T398 T398_D In_12 T356_D VDD pmos w=54.0n l=20n nfin=2 
T400 T400_D In_12 T358_D VDD pmos w=54.0n l=20n nfin=2 
T402 T402_D In_12 T360_D VDD pmos w=54.0n l=20n nfin=2 
T404 T404_D In_12 T362_D VDD pmos w=54.0n l=20n nfin=2 
T406 T406_D In_12 T364_D VDD pmos w=54.0n l=20n nfin=2 
T408 T408_D In_12 T366_D VDD pmos w=54.0n l=20n nfin=2 
T410 T410_D In_12 T368_D VDD pmos w=54.0n l=20n nfin=2 
T412 T412_D In_12 T370_D VDD pmos w=54.0n l=20n nfin=2 
T414 T414_D In_12 T372_D VDD pmos w=54.0n l=20n nfin=2 
T416 T416_D In_12 T374_D VDD pmos w=54.0n l=20n nfin=2 
T418 T418_D In_12 T376_D VDD pmos w=54.0n l=20n nfin=2 
T420 T420_D In_12 T378_D VDD pmos w=54.0n l=20n nfin=2 
T422 T422_D In_12 T380_D VDD pmos w=54.0n l=20n nfin=2 
T424 T424_D In_12 T382_D VDD pmos w=54.0n l=20n nfin=2 
T426 T426_D In_10 T384_D VDD pmos w=54.0n l=20n nfin=2 
T428 T428_D In_10 T386_D VDD pmos w=54.0n l=20n nfin=2 
T430 T430_D In_10 VSS VDD pmos w=54.0n l=20n nfin=2 
T432 T432_D In_10 VSS VDD pmos w=54.0n l=20n nfin=2 
T434 T434_D In_10 VSS VDD pmos w=54.0n l=20n nfin=2 
T436 T436_D In_10 T394_D VDD pmos w=54.0n l=20n nfin=2 
T438 T438_D In_10 T398_D VDD pmos w=54.0n l=20n nfin=2 
T440 T440_D In_10 T402_D VDD pmos w=54.0n l=20n nfin=2 
T442 T442_D In_10 T406_D VDD pmos w=54.0n l=20n nfin=2 
T444 T444_D In_10 T410_D VDD pmos w=54.0n l=20n nfin=2 
T446 T446_D In_10 T414_D VDD pmos w=54.0n l=20n nfin=2 
T448 T448_D In_10 T418_D VDD pmos w=54.0n l=20n nfin=2 
T450 T450_D In_10 T384_D VDD pmos w=54.0n l=20n nfin=2 
T452 T452_D In_10 T386_D VDD pmos w=54.0n l=20n nfin=2 
T454 T454_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T456 T456_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T458 T458_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T460 T460_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T462 T462_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T464 T464_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T466 T466_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T468 T468_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T470 T470_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T472 T472_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T474 T474_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T476 T476_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T478 T478_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T480 T480_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T482 T482_D In_11 VSS VDD pmos w=54.0n l=20n nfin=2 
T484 Y_0 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T486 Y_1 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T488 Y_2 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T490 Y_3 In_1 VDD VDD pmos w=54.0n l=20n nfin=2 
T492 Y_4 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T494 Y_5 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T496 Y_6 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T498 Y_7 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T500 Y_8 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T502 Y_9 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T504 Y_10 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T506 Y_11 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T508 Y_12 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T510 Y_13 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T512 Y_14 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
T514 Y_15 In_1 VSS VDD pmos w=54.0n l=20n nfin=2 
.ENDS

