.SUBCKT xor3_1 In_0 In_1 In_2 VDD VSS Y_0
T1 T0_D In_2 VDD VSS nmos w=54.0n l=20n nfin=2 
T3 T2_D In_2 VSS VSS nmos w=54.0n l=20n nfin=2 
T5 T4_D In_1 T2_D VSS nmos w=54.0n l=20n nfin=2 
T7 T6_D In_1 T0_D VSS nmos w=54.0n l=20n nfin=2 
T9 Y_0 In_0 T6_D VSS nmos w=54.0n l=20n nfin=2 
T0 T0_D In_2 VSS VDD pmos w=54.0n l=20n nfin=2 
T2 T2_D In_2 VDD VDD pmos w=54.0n l=20n nfin=2 
T4 T4_D In_1 T0_D VDD pmos w=54.0n l=20n nfin=2 
T6 T6_D In_1 T2_D VDD pmos w=54.0n l=20n nfin=2 
T8 Y_0 In_0 T4_D VDD pmos w=54.0n l=20n nfin=2 
.ENDS

