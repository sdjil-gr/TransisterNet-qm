.SUBCKT int2float In_0 In_1 In_10 In_2 In_3 In_4 In_5 In_6 In_7 In_8 In_9 VDD VSS Y_0 Y_1 Y_2 Y_3 Y_4 Y_5 Y_6
T1 T0_D In_0 VSS VSS nmos w=54.0n l=20n nfin=2 
T3 T2_D In_4 T0_D VSS nmos w=54.0n l=20n nfin=2 
T5 T4_D In_4 VDD VSS nmos w=54.0n l=20n nfin=2 
T7 T6_D In_4 T0_D VSS nmos w=54.0n l=20n nfin=2 
T9 T8_D In_4 T0_D VSS nmos w=54.0n l=20n nfin=2 
T11 T10_D In_2 T2_D VSS nmos w=54.0n l=20n nfin=2 
T13 T12_D In_2 T4_D VSS nmos w=54.0n l=20n nfin=2 
T15 T14_D In_2 T4_D VSS nmos w=54.0n l=20n nfin=2 
T17 T16_D In_2 T6_D VSS nmos w=54.0n l=20n nfin=2 
T19 T18_D In_2 T6_D VSS nmos w=54.0n l=20n nfin=2 
T21 T20_D In_2 VDD VSS nmos w=54.0n l=20n nfin=2 
T23 T22_D In_2 T6_D VSS nmos w=54.0n l=20n nfin=2 
T25 T24_D In_2 T4_D VSS nmos w=54.0n l=20n nfin=2 
T27 T26_D In_2 T8_D VSS nmos w=54.0n l=20n nfin=2 
T29 T28_D In_3 T10_D VSS nmos w=54.0n l=20n nfin=2 
T31 T30_D In_3 T12_D VSS nmos w=54.0n l=20n nfin=2 
T33 T32_D In_3 T14_D VSS nmos w=54.0n l=20n nfin=2 
T35 T34_D In_3 T14_D VSS nmos w=54.0n l=20n nfin=2 
T37 T36_D In_3 VSS VSS nmos w=54.0n l=20n nfin=2 
T39 T38_D In_3 T16_D VSS nmos w=54.0n l=20n nfin=2 
T41 T40_D In_3 T18_D VSS nmos w=54.0n l=20n nfin=2 
T43 T42_D In_3 T20_D VSS nmos w=54.0n l=20n nfin=2 
T45 T44_D In_3 T14_D VSS nmos w=54.0n l=20n nfin=2 
T47 T46_D In_3 T20_D VSS nmos w=54.0n l=20n nfin=2 
T49 T48_D In_3 T22_D VSS nmos w=54.0n l=20n nfin=2 
T51 T50_D In_3 T24_D VSS nmos w=54.0n l=20n nfin=2 
T53 T52_D In_3 VDD VSS nmos w=54.0n l=20n nfin=2 
T55 T54_D In_3 T26_D VSS nmos w=54.0n l=20n nfin=2 
T57 T56_D In_5 T28_D VSS nmos w=54.0n l=20n nfin=2 
T59 T58_D In_5 T30_D VSS nmos w=54.0n l=20n nfin=2 
T61 T60_D In_5 T32_D VSS nmos w=54.0n l=20n nfin=2 
T63 T62_D In_5 T34_D VSS nmos w=54.0n l=20n nfin=2 
T65 T64_D In_5 T36_D VSS nmos w=54.0n l=20n nfin=2 
T67 T66_D In_5 T28_D VSS nmos w=54.0n l=20n nfin=2 
T69 T68_D In_5 T40_D VSS nmos w=54.0n l=20n nfin=2 
T71 T70_D In_5 T42_D VSS nmos w=54.0n l=20n nfin=2 
T73 T72_D In_5 T34_D VSS nmos w=54.0n l=20n nfin=2 
T75 T74_D In_5 VDD VSS nmos w=54.0n l=20n nfin=2 
T77 T76_D In_5 T44_D VSS nmos w=54.0n l=20n nfin=2 
T79 T78_D In_5 T48_D VSS nmos w=54.0n l=20n nfin=2 
T81 T80_D In_5 T50_D VSS nmos w=54.0n l=20n nfin=2 
T83 T82_D In_5 T32_D VSS nmos w=54.0n l=20n nfin=2 
T85 T84_D In_5 T54_D VSS nmos w=54.0n l=20n nfin=2 
T87 T86_D In_5 T30_D VSS nmos w=54.0n l=20n nfin=2 
T89 T88_D In_5 VDD VSS nmos w=54.0n l=20n nfin=2 
T91 T90_D In_5 T36_D VSS nmos w=54.0n l=20n nfin=2 
T93 T92_D In_6 T58_D VSS nmos w=54.0n l=20n nfin=2 
T95 T94_D In_6 T60_D VSS nmos w=54.0n l=20n nfin=2 
T97 T96_D In_6 T62_D VSS nmos w=54.0n l=20n nfin=2 
T99 T98_D In_6 T64_D VSS nmos w=54.0n l=20n nfin=2 
T101 T100_D In_6 VDD VSS nmos w=54.0n l=20n nfin=2 
T103 T102_D In_6 VDD VSS nmos w=54.0n l=20n nfin=2 
T105 T104_D In_6 T70_D VSS nmos w=54.0n l=20n nfin=2 
T107 T106_D In_6 T72_D VSS nmos w=54.0n l=20n nfin=2 
T109 T108_D In_6 T74_D VSS nmos w=54.0n l=20n nfin=2 
T111 T110_D In_6 T76_D VSS nmos w=54.0n l=20n nfin=2 
T113 T112_D In_6 T80_D VSS nmos w=54.0n l=20n nfin=2 
T115 T114_D In_6 T62_D VSS nmos w=54.0n l=20n nfin=2 
T117 T116_D In_6 T74_D VSS nmos w=54.0n l=20n nfin=2 
T119 T118_D In_6 T82_D VSS nmos w=54.0n l=20n nfin=2 
T121 T120_D In_6 T86_D VSS nmos w=54.0n l=20n nfin=2 
T123 T122_D In_6 T60_D VSS nmos w=54.0n l=20n nfin=2 
T125 T124_D In_6 VDD VSS nmos w=54.0n l=20n nfin=2 
T127 T126_D In_6 T90_D VSS nmos w=54.0n l=20n nfin=2 
T129 T128_D In_8 VSS VSS nmos w=54.0n l=20n nfin=2 
T131 T130_D In_8 T96_D VSS nmos w=54.0n l=20n nfin=2 
T133 T132_D In_8 T98_D VSS nmos w=54.0n l=20n nfin=2 
T135 T134_D In_8 T100_D VSS nmos w=54.0n l=20n nfin=2 
T137 T136_D In_8 VSS VSS nmos w=54.0n l=20n nfin=2 
T139 T138_D In_8 VSS VSS nmos w=54.0n l=20n nfin=2 
T141 T140_D In_8 VDD VSS nmos w=54.0n l=20n nfin=2 
T143 T142_D In_8 T106_D VSS nmos w=54.0n l=20n nfin=2 
T145 T144_D In_8 T108_D VSS nmos w=54.0n l=20n nfin=2 
T147 T146_D In_8 T106_D VSS nmos w=54.0n l=20n nfin=2 
T149 T148_D In_8 T100_D VSS nmos w=54.0n l=20n nfin=2 
T151 T150_D In_8 T114_D VSS nmos w=54.0n l=20n nfin=2 
T153 T152_D In_8 T116_D VSS nmos w=54.0n l=20n nfin=2 
T155 T154_D In_8 T114_D VSS nmos w=54.0n l=20n nfin=2 
T157 T156_D In_8 T100_D VSS nmos w=54.0n l=20n nfin=2 
T159 T158_D In_8 T96_D VSS nmos w=54.0n l=20n nfin=2 
T161 T160_D In_8 T96_D VSS nmos w=54.0n l=20n nfin=2 
T163 T162_D In_8 T116_D VSS nmos w=54.0n l=20n nfin=2 
T165 T164_D In_8 VDD VSS nmos w=54.0n l=20n nfin=2 
T167 T166_D In_8 T126_D VSS nmos w=54.0n l=20n nfin=2 
T169 T168_D In_9 VDD VSS nmos w=54.0n l=20n nfin=2 
T171 T170_D In_9 T132_D VSS nmos w=54.0n l=20n nfin=2 
T173 T172_D In_9 T134_D VSS nmos w=54.0n l=20n nfin=2 
T175 T174_D In_9 VSS VSS nmos w=54.0n l=20n nfin=2 
T177 T176_D In_9 T132_D VSS nmos w=54.0n l=20n nfin=2 
T179 T178_D In_9 VDD VSS nmos w=54.0n l=20n nfin=2 
T181 T180_D In_9 VDD VSS nmos w=54.0n l=20n nfin=2 
T183 T182_D In_9 T144_D VSS nmos w=54.0n l=20n nfin=2 
T185 T184_D In_9 T144_D VSS nmos w=54.0n l=20n nfin=2 
T187 T186_D In_9 T148_D VSS nmos w=54.0n l=20n nfin=2 
T189 T188_D In_9 T140_D VSS nmos w=54.0n l=20n nfin=2 
T191 T190_D In_9 VDD VSS nmos w=54.0n l=20n nfin=2 
T193 T192_D In_9 T152_D VSS nmos w=54.0n l=20n nfin=2 
T195 T194_D In_9 T152_D VSS nmos w=54.0n l=20n nfin=2 
T197 T196_D In_9 T156_D VSS nmos w=54.0n l=20n nfin=2 
T199 T198_D In_9 VDD VSS nmos w=54.0n l=20n nfin=2 
T201 T200_D In_9 T140_D VSS nmos w=54.0n l=20n nfin=2 
T203 T202_D In_9 T140_D VSS nmos w=54.0n l=20n nfin=2 
T205 T204_D In_9 T162_D VSS nmos w=54.0n l=20n nfin=2 
T207 T206_D In_9 T134_D VSS nmos w=54.0n l=20n nfin=2 
T209 T208_D In_9 T140_D VSS nmos w=54.0n l=20n nfin=2 
T211 T210_D In_9 VDD VSS nmos w=54.0n l=20n nfin=2 
T213 T212_D In_9 T166_D VSS nmos w=54.0n l=20n nfin=2 
T215 T214_D In_7 T170_D VSS nmos w=54.0n l=20n nfin=2 
T217 T216_D In_7 T172_D VSS nmos w=54.0n l=20n nfin=2 
T219 T218_D In_7 T176_D VSS nmos w=54.0n l=20n nfin=2 
T221 T220_D In_7 T180_D VSS nmos w=54.0n l=20n nfin=2 
T223 T222_D In_7 T184_D VSS nmos w=54.0n l=20n nfin=2 
T225 T224_D In_7 T186_D VSS nmos w=54.0n l=20n nfin=2 
T227 T226_D In_7 T188_D VSS nmos w=54.0n l=20n nfin=2 
T229 T228_D In_7 T190_D VSS nmos w=54.0n l=20n nfin=2 
T231 T230_D In_7 T194_D VSS nmos w=54.0n l=20n nfin=2 
T233 T232_D In_7 T196_D VSS nmos w=54.0n l=20n nfin=2 
T235 T234_D In_7 T200_D VSS nmos w=54.0n l=20n nfin=2 
T237 T236_D In_7 T178_D VSS nmos w=54.0n l=20n nfin=2 
T239 T238_D In_7 T204_D VSS nmos w=54.0n l=20n nfin=2 
T241 T240_D In_7 T206_D VSS nmos w=54.0n l=20n nfin=2 
T243 T242_D In_7 T208_D VSS nmos w=54.0n l=20n nfin=2 
T245 T244_D In_7 T212_D VSS nmos w=54.0n l=20n nfin=2 
T247 T246_D In_10 T216_D VSS nmos w=54.0n l=20n nfin=2 
T249 T248_D In_10 VDD VSS nmos w=54.0n l=20n nfin=2 
T251 T250_D In_10 VDD VSS nmos w=54.0n l=20n nfin=2 
T253 T252_D In_10 T224_D VSS nmos w=54.0n l=20n nfin=2 
T255 T254_D In_10 T228_D VSS nmos w=54.0n l=20n nfin=2 
T257 T256_D In_10 T232_D VSS nmos w=54.0n l=20n nfin=2 
T259 T258_D In_10 T236_D VSS nmos w=54.0n l=20n nfin=2 
T261 T260_D In_10 T240_D VSS nmos w=54.0n l=20n nfin=2 
T263 T262_D In_10 VDD VSS nmos w=54.0n l=20n nfin=2 
T265 T264_D In_10 VDD VSS nmos w=54.0n l=20n nfin=2 
T267 Y_0 In_1 VDD VSS nmos w=54.0n l=20n nfin=2 
T269 Y_1 In_1 VDD VSS nmos w=54.0n l=20n nfin=2 
T271 Y_2 In_1 VDD VSS nmos w=54.0n l=20n nfin=2 
T273 Y_3 In_1 T254_D VSS nmos w=54.0n l=20n nfin=2 
T275 Y_4 In_1 T258_D VSS nmos w=54.0n l=20n nfin=2 
T277 Y_5 In_1 T262_D VSS nmos w=54.0n l=20n nfin=2 
T279 Y_6 In_1 VDD VSS nmos w=54.0n l=20n nfin=2 
T0 T0_D In_0 VSS VDD pmos w=54.0n l=20n nfin=2 
T2 T2_D In_4 VDD VDD pmos w=54.0n l=20n nfin=2 
T4 T4_D In_4 VSS VDD pmos w=54.0n l=20n nfin=2 
T6 T6_D In_4 T0_D VDD pmos w=54.0n l=20n nfin=2 
T8 T8_D In_4 T0_D VDD pmos w=54.0n l=20n nfin=2 
T10 T10_D In_2 VDD VDD pmos w=54.0n l=20n nfin=2 
T12 T12_D In_2 VSS VDD pmos w=54.0n l=20n nfin=2 
T14 T14_D In_2 T4_D VDD pmos w=54.0n l=20n nfin=2 
T16 T16_D In_2 T6_D VDD pmos w=54.0n l=20n nfin=2 
T18 T18_D In_2 T6_D VDD pmos w=54.0n l=20n nfin=2 
T20 T20_D In_2 VSS VDD pmos w=54.0n l=20n nfin=2 
T22 T22_D In_2 VSS VDD pmos w=54.0n l=20n nfin=2 
T24 T24_D In_2 T4_D VDD pmos w=54.0n l=20n nfin=2 
T26 T26_D In_2 T4_D VDD pmos w=54.0n l=20n nfin=2 
T28 T28_D In_3 VDD VDD pmos w=54.0n l=20n nfin=2 
T30 T30_D In_3 VSS VDD pmos w=54.0n l=20n nfin=2 
T32 T32_D In_3 VDD VDD pmos w=54.0n l=20n nfin=2 
T34 T34_D In_3 T14_D VDD pmos w=54.0n l=20n nfin=2 
T36 T36_D In_3 T14_D VDD pmos w=54.0n l=20n nfin=2 
T38 T38_D In_3 T16_D VDD pmos w=54.0n l=20n nfin=2 
T40 T40_D In_3 T18_D VDD pmos w=54.0n l=20n nfin=2 
T42 T42_D In_3 T20_D VDD pmos w=54.0n l=20n nfin=2 
T44 T44_D In_3 T14_D VDD pmos w=54.0n l=20n nfin=2 
T46 T46_D In_3 T20_D VDD pmos w=54.0n l=20n nfin=2 
T48 T48_D In_3 T22_D VDD pmos w=54.0n l=20n nfin=2 
T50 T50_D In_3 T14_D VDD pmos w=54.0n l=20n nfin=2 
T52 T52_D In_3 VSS VDD pmos w=54.0n l=20n nfin=2 
T54 T54_D In_3 T14_D VDD pmos w=54.0n l=20n nfin=2 
T56 T56_D In_5 VSS VDD pmos w=54.0n l=20n nfin=2 
T58 T58_D In_5 VSS VDD pmos w=54.0n l=20n nfin=2 
T60 T60_D In_5 VDD VDD pmos w=54.0n l=20n nfin=2 
T62 T62_D In_5 VSS VDD pmos w=54.0n l=20n nfin=2 
T64 T64_D In_5 VDD VDD pmos w=54.0n l=20n nfin=2 
T66 T66_D In_5 VSS VDD pmos w=54.0n l=20n nfin=2 
T68 T68_D In_5 T38_D VDD pmos w=54.0n l=20n nfin=2 
T70 T70_D In_5 T42_D VDD pmos w=54.0n l=20n nfin=2 
T72 T72_D In_5 T34_D VDD pmos w=54.0n l=20n nfin=2 
T74 T74_D In_5 VSS VDD pmos w=54.0n l=20n nfin=2 
T76 T76_D In_5 T44_D VDD pmos w=54.0n l=20n nfin=2 
T78 T78_D In_5 T46_D VDD pmos w=54.0n l=20n nfin=2 
T80 T80_D In_5 T50_D VDD pmos w=54.0n l=20n nfin=2 
T82 T82_D In_5 T32_D VDD pmos w=54.0n l=20n nfin=2 
T84 T84_D In_5 T52_D VDD pmos w=54.0n l=20n nfin=2 
T86 T86_D In_5 T30_D VDD pmos w=54.0n l=20n nfin=2 
T88 T88_D In_5 T34_D VDD pmos w=54.0n l=20n nfin=2 
T90 T90_D In_5 VDD VDD pmos w=54.0n l=20n nfin=2 
T92 T92_D In_6 T56_D VDD pmos w=54.0n l=20n nfin=2 
T94 T94_D In_6 VDD VDD pmos w=54.0n l=20n nfin=2 
T96 T96_D In_6 VSS VDD pmos w=54.0n l=20n nfin=2 
T98 T98_D In_6 VDD VDD pmos w=54.0n l=20n nfin=2 
T100 T100_D In_6 VSS VDD pmos w=54.0n l=20n nfin=2 
T102 T102_D In_6 T66_D VDD pmos w=54.0n l=20n nfin=2 
T104 T104_D In_6 T68_D VDD pmos w=54.0n l=20n nfin=2 
T106 T106_D In_6 T72_D VDD pmos w=54.0n l=20n nfin=2 
T108 T108_D In_6 T74_D VDD pmos w=54.0n l=20n nfin=2 
T110 T110_D In_6 T76_D VDD pmos w=54.0n l=20n nfin=2 
T112 T112_D In_6 T78_D VDD pmos w=54.0n l=20n nfin=2 
T114 T114_D In_6 T62_D VDD pmos w=54.0n l=20n nfin=2 
T116 T116_D In_6 VSS VDD pmos w=54.0n l=20n nfin=2 
T118 T118_D In_6 T82_D VDD pmos w=54.0n l=20n nfin=2 
T120 T120_D In_6 T84_D VDD pmos w=54.0n l=20n nfin=2 
T122 T122_D In_6 T60_D VDD pmos w=54.0n l=20n nfin=2 
T124 T124_D In_6 T88_D VDD pmos w=54.0n l=20n nfin=2 
T126 T126_D In_6 VDD VDD pmos w=54.0n l=20n nfin=2 
T128 T128_D In_8 T92_D VDD pmos w=54.0n l=20n nfin=2 
T130 T130_D In_8 T94_D VDD pmos w=54.0n l=20n nfin=2 
T132 T132_D In_8 VDD VDD pmos w=54.0n l=20n nfin=2 
T134 T134_D In_8 VSS VDD pmos w=54.0n l=20n nfin=2 
T136 T136_D In_8 T102_D VDD pmos w=54.0n l=20n nfin=2 
T138 T138_D In_8 T94_D VDD pmos w=54.0n l=20n nfin=2 
T140 T140_D In_8 VSS VDD pmos w=54.0n l=20n nfin=2 
T142 T142_D In_8 T104_D VDD pmos w=54.0n l=20n nfin=2 
T144 T144_D In_8 T108_D VDD pmos w=54.0n l=20n nfin=2 
T146 T146_D In_8 T110_D VDD pmos w=54.0n l=20n nfin=2 
T148 T148_D In_8 T100_D VDD pmos w=54.0n l=20n nfin=2 
T150 T150_D In_8 T112_D VDD pmos w=54.0n l=20n nfin=2 
T152 T152_D In_8 T116_D VDD pmos w=54.0n l=20n nfin=2 
T154 T154_D In_8 T118_D VDD pmos w=54.0n l=20n nfin=2 
T156 T156_D In_8 T100_D VDD pmos w=54.0n l=20n nfin=2 
T158 T158_D In_8 T120_D VDD pmos w=54.0n l=20n nfin=2 
T160 T160_D In_8 T122_D VDD pmos w=54.0n l=20n nfin=2 
T162 T162_D In_8 T116_D VDD pmos w=54.0n l=20n nfin=2 
T164 T164_D In_8 T124_D VDD pmos w=54.0n l=20n nfin=2 
T166 T166_D In_8 VDD VDD pmos w=54.0n l=20n nfin=2 
T168 T168_D In_9 T128_D VDD pmos w=54.0n l=20n nfin=2 
T170 T170_D In_9 T130_D VDD pmos w=54.0n l=20n nfin=2 
T172 T172_D In_9 VSS VDD pmos w=54.0n l=20n nfin=2 
T174 T174_D In_9 T136_D VDD pmos w=54.0n l=20n nfin=2 
T176 T176_D In_9 T138_D VDD pmos w=54.0n l=20n nfin=2 
T178 T178_D In_9 T140_D VDD pmos w=54.0n l=20n nfin=2 
T180 T180_D In_9 T138_D VDD pmos w=54.0n l=20n nfin=2 
T182 T182_D In_9 T142_D VDD pmos w=54.0n l=20n nfin=2 
T184 T184_D In_9 T146_D VDD pmos w=54.0n l=20n nfin=2 
T186 T186_D In_9 T148_D VDD pmos w=54.0n l=20n nfin=2 
T188 T188_D In_9 T140_D VDD pmos w=54.0n l=20n nfin=2 
T190 T190_D In_9 T140_D VDD pmos w=54.0n l=20n nfin=2 
T192 T192_D In_9 T150_D VDD pmos w=54.0n l=20n nfin=2 
T194 T194_D In_9 T154_D VDD pmos w=54.0n l=20n nfin=2 
T196 T196_D In_9 T156_D VDD pmos w=54.0n l=20n nfin=2 
T198 T198_D In_9 VSS VDD pmos w=54.0n l=20n nfin=2 
T200 T200_D In_9 T140_D VDD pmos w=54.0n l=20n nfin=2 
T202 T202_D In_9 T158_D VDD pmos w=54.0n l=20n nfin=2 
T204 T204_D In_9 T160_D VDD pmos w=54.0n l=20n nfin=2 
T206 T206_D In_9 T134_D VDD pmos w=54.0n l=20n nfin=2 
T208 T208_D In_9 VSS VDD pmos w=54.0n l=20n nfin=2 
T210 T210_D In_9 T164_D VDD pmos w=54.0n l=20n nfin=2 
T212 T212_D In_9 VDD VDD pmos w=54.0n l=20n nfin=2 
T214 T214_D In_7 T168_D VDD pmos w=54.0n l=20n nfin=2 
T216 T216_D In_7 VSS VDD pmos w=54.0n l=20n nfin=2 
T218 T218_D In_7 T174_D VDD pmos w=54.0n l=20n nfin=2 
T220 T220_D In_7 T178_D VDD pmos w=54.0n l=20n nfin=2 
T222 T222_D In_7 T182_D VDD pmos w=54.0n l=20n nfin=2 
T224 T224_D In_7 T186_D VDD pmos w=54.0n l=20n nfin=2 
T226 T226_D In_7 T188_D VDD pmos w=54.0n l=20n nfin=2 
T228 T228_D In_7 T188_D VDD pmos w=54.0n l=20n nfin=2 
T230 T230_D In_7 T192_D VDD pmos w=54.0n l=20n nfin=2 
T232 T232_D In_7 T188_D VDD pmos w=54.0n l=20n nfin=2 
T234 T234_D In_7 T198_D VDD pmos w=54.0n l=20n nfin=2 
T236 T236_D In_7 T198_D VDD pmos w=54.0n l=20n nfin=2 
T238 T238_D In_7 T202_D VDD pmos w=54.0n l=20n nfin=2 
T240 T240_D In_7 T198_D VDD pmos w=54.0n l=20n nfin=2 
T242 T242_D In_7 VSS VDD pmos w=54.0n l=20n nfin=2 
T244 T244_D In_7 T210_D VDD pmos w=54.0n l=20n nfin=2 
T246 T246_D In_10 T214_D VDD pmos w=54.0n l=20n nfin=2 
T248 T248_D In_10 T218_D VDD pmos w=54.0n l=20n nfin=2 
T250 T250_D In_10 T220_D VDD pmos w=54.0n l=20n nfin=2 
T252 T252_D In_10 T222_D VDD pmos w=54.0n l=20n nfin=2 
T254 T254_D In_10 T226_D VDD pmos w=54.0n l=20n nfin=2 
T256 T256_D In_10 T230_D VDD pmos w=54.0n l=20n nfin=2 
T258 T258_D In_10 T234_D VDD pmos w=54.0n l=20n nfin=2 
T260 T260_D In_10 T238_D VDD pmos w=54.0n l=20n nfin=2 
T262 T262_D In_10 T242_D VDD pmos w=54.0n l=20n nfin=2 
T264 T264_D In_10 T244_D VDD pmos w=54.0n l=20n nfin=2 
T266 Y_0 In_1 T246_D VDD pmos w=54.0n l=20n nfin=2 
T268 Y_1 In_1 T248_D VDD pmos w=54.0n l=20n nfin=2 
T270 Y_2 In_1 T250_D VDD pmos w=54.0n l=20n nfin=2 
T272 Y_3 In_1 T252_D VDD pmos w=54.0n l=20n nfin=2 
T274 Y_4 In_1 T256_D VDD pmos w=54.0n l=20n nfin=2 
T276 Y_5 In_1 T260_D VDD pmos w=54.0n l=20n nfin=2 
T278 Y_6 In_1 T264_D VDD pmos w=54.0n l=20n nfin=2 
.ENDS

